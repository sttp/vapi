module version

const (
	sttpsource     = 'STTP V Library'
	sttpversion    = '0.0.1'
	sttpupdated_on = '2023-04-19'
)
