module parser
import encoding
import github.com.antlr.antlr4.runtime.Go.antlr
const (
_=fmt.printf 
_=unicode.is_letter 
serialized_lexer_atn=[u16(3 ,) ,24715 ,42794 ,33075 ,47597 ,16764 ,15335 ,30598 ,22884 ,2 ,100 ,992 ,8 ,1 ,4 ,2 ,9 ,2 ,4 ,3 ,9 ,3 ,4 ,4 ,9 ,4 ,4 ,5 ,9 ,5 ,4 ,6 ,9 ,6 ,4 ,7 ,9 ,7 ,4 ,8 ,9 ,8 ,4 ,9 ,9 ,9 ,4 ,10 ,9 ,10 ,4 ,11 ,9 ,11 ,4 ,12 ,9 ,12 ,4 ,13 ,9 ,13 ,4 ,14 ,9 ,14 ,4 ,15 ,9 ,15 ,4 ,16 ,9 ,16 ,4 ,17 ,9 ,17 ,4 ,18 ,9 ,18 ,4 ,19 ,9 ,19 ,4 ,20 ,9 ,20 ,4 ,21 ,9 ,21 ,4 ,22 ,9 ,22 ,4 ,23 ,9 ,23 ,4 ,24 ,9 ,24 ,4 ,25 ,9 ,25 ,4 ,26 ,9 ,26 ,4 ,27 ,9 ,27 ,4 ,28 ,9 ,28 ,4 ,29 ,9 ,29 ,4 ,30 ,9 ,30 ,4 ,31 ,9 ,31 ,4 ,32 ,9 ,32 ,4 ,33 ,9 ,33 ,4 ,34 ,9 ,34 ,4 ,35 ,9 ,35 ,4 ,36 ,9 ,36 ,4 ,37 ,9 ,37 ,4 ,38 ,9 ,38 ,4 ,39 ,9 ,39 ,4 ,40 ,9 ,40 ,4 ,41 ,9 ,41 ,4 ,42 ,9 ,42 ,4 ,43 ,9 ,43 ,4 ,44 ,9 ,44 ,4 ,45 ,9 ,45 ,4 ,46 ,9 ,46 ,4 ,47 ,9 ,47 ,4 ,48 ,9 ,48 ,4 ,49 ,9 ,49 ,4 ,50 ,9 ,50 ,4 ,51 ,9 ,51 ,4 ,52 ,9 ,52 ,4 ,53 ,9 ,53 ,4 ,54 ,9 ,54 ,4 ,55 ,9 ,55 ,4 ,56 ,9 ,56 ,4 ,57 ,9 ,57 ,4 ,58 ,9 ,58 ,4 ,59 ,9 ,59 ,4 ,60 ,9 ,60 ,4 ,61 ,9 ,61 ,4 ,62 ,9 ,62 ,4 ,63 ,9 ,63 ,4 ,64 ,9 ,64 ,4 ,65 ,9 ,65 ,4 ,66 ,9 ,66 ,4 ,67 ,9 ,67 ,4 ,68 ,9 ,68 ,4 ,69 ,9 ,69 ,4 ,70 ,9 ,70 ,4 ,71 ,9 ,71 ,4 ,72 ,9 ,72 ,4 ,73 ,9 ,73 ,4 ,74 ,9 ,74 ,4 ,75 ,9 ,75 ,4 ,76 ,9 ,76 ,4 ,77 ,9 ,77 ,4 ,78 ,9 ,78 ,4 ,79 ,9 ,79 ,4 ,80 ,9 ,80 ,4 ,81 ,9 ,81 ,4 ,82 ,9 ,82 ,4 ,83 ,9 ,83 ,4 ,84 ,9 ,84 ,4 ,85 ,9 ,85 ,4 ,86 ,9 ,86 ,4 ,87 ,9 ,87 ,4 ,88 ,9 ,88 ,4 ,89 ,9 ,89 ,4 ,90 ,9 ,90 ,4 ,91 ,9 ,91 ,4 ,92 ,9 ,92 ,4 ,93 ,9 ,93 ,4 ,94 ,9 ,94 ,4 ,95 ,9 ,95 ,4 ,96 ,9 ,96 ,4 ,97 ,9 ,97 ,4 ,98 ,9 ,98 ,4 ,99 ,9 ,99 ,4 ,100 ,9 ,100 ,4 ,101 ,9 ,101 ,4 ,102 ,9 ,102 ,4 ,103 ,9 ,103 ,4 ,104 ,9 ,104 ,4 ,105 ,9 ,105 ,4 ,106 ,9 ,106 ,4 ,107 ,9 ,107 ,4 ,108 ,9 ,108 ,4 ,109 ,9 ,109 ,4 ,110 ,9 ,110 ,4 ,111 ,9 ,111 ,4 ,112 ,9 ,112 ,4 ,113 ,9 ,113 ,4 ,114 ,9 ,114 ,4 ,115 ,9 ,115 ,4 ,116 ,9 ,116 ,4 ,117 ,9 ,117 ,4 ,118 ,9 ,118 ,4 ,119 ,9 ,119 ,4 ,120 ,9 ,120 ,4 ,121 ,9 ,121 ,4 ,122 ,9 ,122 ,4 ,123 ,9 ,123 ,4 ,124 ,9 ,124 ,4 ,125 ,9 ,125 ,4 ,126 ,9 ,126 ,4 ,127 ,9 ,127 ,4 ,128 ,9 ,128 ,4 ,129 ,9 ,129 ,3 ,2 ,3 ,2 ,3 ,3 ,3 ,3 ,3 ,4 ,3 ,4 ,3 ,5 ,3 ,5 ,3 ,6 ,3 ,6 ,3 ,7 ,3 ,7 ,3 ,8 ,3 ,8 ,3 ,9 ,3 ,9 ,3 ,10 ,3 ,10 ,3 ,10 ,3 ,10 ,3 ,11 ,3 ,11 ,3 ,12 ,3 ,12 ,3 ,12 ,3 ,13 ,3 ,13 ,3 ,14 ,3 ,14 ,3 ,14 ,3 ,15 ,3 ,15 ,3 ,16 ,3 ,16 ,3 ,16 ,3 ,17 ,3 ,17 ,3 ,17 ,3 ,18 ,3 ,18 ,3 ,18 ,3 ,18 ,3 ,19 ,3 ,19 ,3 ,19 ,3 ,20 ,3 ,20 ,3 ,20 ,3 ,21 ,3 ,21 ,3 ,21 ,3 ,22 ,3 ,22 ,3 ,22 ,3 ,23 ,3 ,23 ,3 ,23 ,3 ,24 ,3 ,24 ,3 ,25 ,3 ,25 ,3 ,26 ,3 ,26 ,3 ,27 ,3 ,27 ,3 ,28 ,3 ,28 ,3 ,29 ,3 ,29 ,3 ,30 ,3 ,30 ,3 ,30 ,3 ,30 ,3 ,31 ,3 ,31 ,3 ,31 ,3 ,31 ,3 ,32 ,3 ,32 ,3 ,32 ,3 ,32 ,3 ,33 ,3 ,33 ,3 ,33 ,3 ,33 ,3 ,33 ,3 ,33 ,3 ,33 ,3 ,34 ,3 ,34 ,3 ,34 ,3 ,35 ,3 ,35 ,3 ,35 ,3 ,35 ,3 ,35 ,3 ,35 ,3 ,35 ,3 ,35 ,3 ,36 ,3 ,36 ,3 ,36 ,3 ,36 ,3 ,36 ,3 ,36 ,3 ,36 ,3 ,36 ,3 ,36 ,3 ,37 ,3 ,37 ,3 ,37 ,3 ,37 ,3 ,37 ,3 ,37 ,3 ,37 ,3 ,37 ,3 ,38 ,3 ,38 ,3 ,38 ,3 ,38 ,3 ,38 ,3 ,38 ,3 ,38 ,3 ,38 ,3 ,38 ,3 ,39 ,3 ,39 ,3 ,39 ,3 ,39 ,3 ,39 ,3 ,39 ,3 ,39 ,3 ,39 ,3 ,40 ,3 ,40 ,3 ,40 ,3 ,40 ,3 ,40 ,3 ,40 ,3 ,40 ,3 ,40 ,3 ,40 ,3 ,41 ,3 ,41 ,3 ,41 ,3 ,41 ,3 ,41 ,3 ,41 ,3 ,41 ,3 ,41 ,3 ,41 ,3 ,42 ,3 ,42 ,3 ,42 ,3 ,42 ,3 ,42 ,3 ,43 ,3 ,43 ,3 ,43 ,3 ,43 ,3 ,43 ,3 ,43 ,3 ,43 ,3 ,43 ,3 ,43 ,3 ,44 ,3 ,44 ,3 ,44 ,3 ,44 ,3 ,44 ,3 ,44 ,3 ,44 ,3 ,45 ,3 ,45 ,3 ,45 ,3 ,45 ,3 ,45 ,3 ,45 ,3 ,46 ,3 ,46 ,3 ,46 ,3 ,46 ,3 ,47 ,3 ,47 ,3 ,47 ,3 ,48 ,3 ,48 ,3 ,48 ,3 ,48 ,3 ,48 ,3 ,48 ,3 ,48 ,3 ,48 ,3 ,49 ,3 ,49 ,3 ,49 ,3 ,50 ,3 ,50 ,3 ,50 ,3 ,50 ,3 ,50 ,3 ,50 ,3 ,50 ,3 ,51 ,3 ,51 ,3 ,51 ,3 ,51 ,3 ,51 ,3 ,51 ,3 ,51 ,3 ,51 ,3 ,51 ,3 ,51 ,3 ,52 ,3 ,52 ,3 ,52 ,3 ,52 ,3 ,52 ,3 ,52 ,3 ,52 ,3 ,53 ,3 ,53 ,3 ,53 ,3 ,53 ,3 ,53 ,3 ,53 ,3 ,53 ,3 ,54 ,3 ,54 ,3 ,54 ,3 ,54 ,3 ,54 ,3 ,54 ,3 ,54 ,3 ,54 ,3 ,54 ,3 ,54 ,3 ,55 ,3 ,55 ,3 ,55 ,3 ,55 ,3 ,55 ,3 ,55 ,3 ,55 ,3 ,55 ,3 ,55 ,3 ,55 ,3 ,55 ,3 ,55 ,3 ,56 ,3 ,56 ,3 ,56 ,3 ,56 ,3 ,57 ,3 ,57 ,3 ,57 ,3 ,57 ,3 ,57 ,3 ,58 ,3 ,58 ,3 ,58 ,3 ,58 ,3 ,58 ,3 ,58 ,3 ,59 ,3 ,59 ,3 ,59 ,3 ,59 ,3 ,59 ,3 ,59 ,3 ,60 ,3 ,60 ,3 ,60 ,3 ,60 ,3 ,60 ,3 ,60 ,3 ,61 ,3 ,61 ,3 ,61 ,3 ,61 ,3 ,62 ,3 ,62 ,3 ,62 ,3 ,62 ,3 ,63 ,3 ,63 ,3 ,63 ,3 ,63 ,3 ,63 ,3 ,63 ,3 ,63 ,3 ,63 ,3 ,63 ,3 ,63 ,3 ,63 ,3 ,64 ,3 ,64 ,3 ,64 ,3 ,64 ,3 ,64 ,3 ,65 ,3 ,65 ,3 ,65 ,3 ,66 ,3 ,66 ,3 ,66 ,3 ,66 ,3 ,66 ,3 ,66 ,3 ,67 ,3 ,67 ,3 ,67 ,3 ,67 ,3 ,67 ,3 ,67 ,3 ,68 ,3 ,68 ,3 ,68 ,3 ,68 ,3 ,68 ,3 ,68 ,3 ,68 ,3 ,68 ,3 ,68 ,3 ,68 ,3 ,68 ,3 ,69 ,3 ,69 ,3 ,69 ,3 ,69 ,3 ,69 ,3 ,69 ,3 ,69 ,3 ,69 ,3 ,69 ,3 ,70 ,3 ,70 ,3 ,70 ,3 ,70 ,3 ,70 ,3 ,70 ,3 ,70 ,3 ,70 ,3 ,71 ,3 ,71 ,3 ,71 ,3 ,71 ,3 ,71 ,3 ,71 ,3 ,71 ,3 ,71 ,3 ,72 ,3 ,72 ,3 ,72 ,3 ,72 ,3 ,72 ,3 ,72 ,3 ,73 ,3 ,73 ,3 ,73 ,3 ,73 ,3 ,73 ,3 ,74 ,3 ,74 ,3 ,74 ,3 ,74 ,3 ,74 ,3 ,74 ,3 ,75 ,3 ,75 ,3 ,75 ,3 ,75 ,3 ,75 ,3 ,75 ,3 ,75 ,3 ,75 ,3 ,75 ,3 ,75 ,3 ,75 ,3 ,76 ,3 ,76 ,3 ,76 ,3 ,76 ,3 ,76 ,3 ,76 ,3 ,76 ,3 ,76 ,3 ,76 ,3 ,77 ,3 ,77 ,3 ,77 ,3 ,77 ,3 ,77 ,3 ,77 ,3 ,77 ,3 ,78 ,3 ,78 ,3 ,78 ,3 ,78 ,3 ,78 ,3 ,78 ,3 ,78 ,3 ,79 ,3 ,79 ,3 ,79 ,3 ,79 ,3 ,80 ,3 ,80 ,3 ,80 ,3 ,80 ,3 ,80 ,3 ,81 ,3 ,81 ,3 ,81 ,3 ,81 ,3 ,81 ,3 ,81 ,3 ,81 ,3 ,81 ,3 ,81 ,3 ,82 ,3 ,82 ,3 ,82 ,3 ,82 ,3 ,82 ,3 ,82 ,3 ,82 ,3 ,82 ,3 ,82 ,3 ,82 ,3 ,83 ,3 ,83 ,3 ,83 ,3 ,83 ,3 ,83 ,3 ,83 ,3 ,84 ,3 ,84 ,3 ,84 ,3 ,84 ,3 ,84 ,3 ,84 ,3 ,84 ,3 ,85 ,3 ,85 ,3 ,85 ,3 ,85 ,3 ,85 ,3 ,85 ,3 ,86 ,3 ,86 ,3 ,86 ,3 ,86 ,3 ,87 ,3 ,87 ,3 ,87 ,3 ,87 ,3 ,87 ,3 ,87 ,3 ,87 ,3 ,87 ,3 ,87 ,3 ,87 ,3 ,87 ,5 ,87 ,724 ,10 ,87 ,3 ,88 ,3 ,88 ,6 ,88 ,728 ,10 ,88 ,13 ,88 ,14 ,88 ,729 ,3 ,88 ,3 ,88 ,3 ,88 ,6 ,88 ,735 ,10 ,88 ,13 ,88 ,14 ,88 ,736 ,3 ,88 ,3 ,88 ,3 ,88 ,7 ,88 ,742 ,10 ,88 ,12 ,88 ,14 ,88 ,745 ,11 ,88 ,5 ,88 ,747 ,10 ,88 ,3 ,89 ,6 ,89 ,750 ,10 ,89 ,13 ,89 ,14 ,89 ,751 ,3 ,89 ,3 ,89 ,3 ,89 ,6 ,89 ,757 ,10 ,89 ,13 ,89 ,14 ,89 ,758 ,5 ,89 ,761 ,10 ,89 ,3 ,90 ,6 ,90 ,764 ,10 ,90 ,13 ,90 ,14 ,90 ,765 ,3 ,90 ,3 ,90 ,7 ,90 ,770 ,10 ,90 ,12 ,90 ,14 ,90 ,773 ,11 ,90 ,5 ,90 ,775 ,10 ,90 ,3 ,90 ,3 ,90 ,5 ,90 ,779 ,10 ,90 ,3 ,90 ,6 ,90 ,782 ,10 ,90 ,13 ,90 ,14 ,90 ,783 ,5 ,90 ,786 ,10 ,90 ,3 ,90 ,3 ,90 ,6 ,90 ,790 ,10 ,90 ,13 ,90 ,14 ,90 ,791 ,3 ,90 ,3 ,90 ,5 ,90 ,796 ,10 ,90 ,3 ,90 ,6 ,90 ,799 ,10 ,90 ,13 ,90 ,14 ,90 ,800 ,5 ,90 ,803 ,10 ,90 ,5 ,90 ,805 ,10 ,90 ,3 ,91 ,3 ,91 ,3 ,91 ,3 ,91 ,3 ,91 ,3 ,91 ,3 ,91 ,3 ,91 ,3 ,91 ,5 ,91 ,816 ,10 ,91 ,3 ,92 ,6 ,92 ,819 ,10 ,92 ,13 ,92 ,14 ,92 ,820 ,3 ,92 ,3 ,92 ,6 ,92 ,825 ,10 ,92 ,13 ,92 ,14 ,92 ,826 ,3 ,93 ,3 ,93 ,6 ,93 ,831 ,10 ,93 ,13 ,93 ,14 ,93 ,832 ,3 ,93 ,3 ,93 ,3 ,94 ,3 ,94 ,3 ,94 ,3 ,94 ,7 ,94 ,841 ,10 ,94 ,12 ,94 ,14 ,94 ,844 ,11 ,94 ,3 ,94 ,3 ,94 ,3 ,95 ,3 ,95 ,6 ,95 ,850 ,10 ,95 ,13 ,95 ,14 ,95 ,851 ,3 ,95 ,3 ,95 ,3 ,96 ,3 ,96 ,3 ,96 ,3 ,96 ,7 ,96 ,860 ,10 ,96 ,12 ,96 ,14 ,96 ,863 ,11 ,96 ,3 ,96 ,3 ,96 ,3 ,97 ,3 ,97 ,3 ,97 ,3 ,97 ,7 ,97 ,871 ,10 ,97 ,12 ,97 ,14 ,97 ,874 ,11 ,97 ,3 ,97 ,3 ,97 ,3 ,97 ,5 ,97 ,879 ,10 ,97 ,3 ,97 ,3 ,97 ,3 ,98 ,3 ,98 ,3 ,98 ,3 ,98 ,3 ,99 ,3 ,99 ,3 ,100 ,3 ,100 ,3 ,101 ,3 ,101 ,3 ,102 ,5 ,102 ,894 ,10 ,102 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,5 ,103 ,905 ,10 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,5 ,103 ,912 ,10 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,5 ,103 ,919 ,10 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,5 ,103 ,926 ,10 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,103 ,3 ,104 ,3 ,104 ,3 ,105 ,3 ,105 ,3 ,106 ,3 ,106 ,3 ,107 ,3 ,107 ,3 ,108 ,3 ,108 ,3 ,109 ,3 ,109 ,3 ,110 ,3 ,110 ,3 ,111 ,3 ,111 ,3 ,112 ,3 ,112 ,3 ,113 ,3 ,113 ,3 ,114 ,3 ,114 ,3 ,115 ,3 ,115 ,3 ,116 ,3 ,116 ,3 ,117 ,3 ,117 ,3 ,118 ,3 ,118 ,3 ,119 ,3 ,119 ,3 ,120 ,3 ,120 ,3 ,121 ,3 ,121 ,3 ,122 ,3 ,122 ,3 ,123 ,3 ,123 ,3 ,124 ,3 ,124 ,3 ,125 ,3 ,125 ,3 ,126 ,3 ,126 ,3 ,127 ,3 ,127 ,3 ,128 ,3 ,128 ,3 ,129 ,3 ,129 ,3 ,872 ,2 ,130 ,3 ,3 ,5 ,4 ,7 ,5 ,9 ,6 ,11 ,7 ,13 ,8 ,15 ,9 ,17 ,10 ,19 ,11 ,21 ,12 ,23 ,13 ,25 ,14 ,27 ,15 ,29 ,16 ,31 ,17 ,33 ,18 ,35 ,19 ,37 ,20 ,39 ,21 ,41 ,22 ,43 ,23 ,45 ,24 ,47 ,25 ,49 ,26 ,51 ,27 ,53 ,28 ,55 ,29 ,57 ,30 ,59 ,31 ,61 ,32 ,63 ,33 ,65 ,34 ,67 ,35 ,69 ,36 ,71 ,37 ,73 ,38 ,75 ,39 ,77 ,40 ,79 ,41 ,81 ,42 ,83 ,43 ,85 ,44 ,87 ,45 ,89 ,46 ,91 ,47 ,93 ,48 ,95 ,49 ,97 ,50 ,99 ,51 ,101 ,52 ,103 ,53 ,105 ,54 ,107 ,55 ,109 ,56 ,111 ,57 ,113 ,58 ,115 ,59 ,117 ,60 ,119 ,61 ,121 ,62 ,123 ,63 ,125 ,64 ,127 ,65 ,129 ,66 ,131 ,67 ,133 ,68 ,135 ,69 ,137 ,70 ,139 ,71 ,141 ,72 ,143 ,73 ,145 ,74 ,147 ,75 ,149 ,76 ,151 ,77 ,153 ,78 ,155 ,79 ,157 ,80 ,159 ,81 ,161 ,82 ,163 ,83 ,165 ,84 ,167 ,85 ,169 ,86 ,171 ,87 ,173 ,88 ,175 ,89 ,177 ,90 ,179 ,91 ,181 ,92 ,183 ,93 ,185 ,94 ,187 ,95 ,189 ,96 ,191 ,97 ,193 ,98 ,195 ,99 ,197 ,100 ,199 ,2 ,201 ,2 ,203 ,2 ,205 ,2 ,207 ,2 ,209 ,2 ,211 ,2 ,213 ,2 ,215 ,2 ,217 ,2 ,219 ,2 ,221 ,2 ,223 ,2 ,225 ,2 ,227 ,2 ,229 ,2 ,231 ,2 ,233 ,2 ,235 ,2 ,237 ,2 ,239 ,2 ,241 ,2 ,243 ,2 ,245 ,2 ,247 ,2 ,249 ,2 ,251 ,2 ,253 ,2 ,255 ,2 ,257 ,2 ,3 ,2 ,40 ,3 ,2 ,98 ,98 ,3 ,2 ,95 ,95 ,5 ,2 ,67 ,92 ,97 ,97 ,99 ,124 ,6 ,2 ,50 ,59 ,67 ,92 ,97 ,97 ,99 ,124 ,4 ,2 ,45 ,45 ,47 ,47 ,3 ,2 ,41 ,41 ,3 ,2 ,37 ,37 ,4 ,2 ,12 ,12 ,15 ,15 ,5 ,2 ,11 ,13 ,15 ,15 ,34 ,34 ,3 ,2 ,50 ,59 ,5 ,2 ,50 ,59 ,67 ,72 ,99 ,104 ,9 ,2 ,35 ,35 ,37 ,38 ,47 ,48 ,50 ,59 ,66 ,92 ,97 ,97 ,99 ,124 ,4 ,2 ,67 ,67 ,99 ,99 ,4 ,2 ,68 ,68 ,100 ,100 ,4 ,2 ,69 ,69 ,101 ,101 ,4 ,2 ,70 ,70 ,102 ,102 ,4 ,2 ,71 ,71 ,103 ,103 ,4 ,2 ,72 ,72 ,104 ,104 ,4 ,2 ,73 ,73 ,105 ,105 ,4 ,2 ,74 ,74 ,106 ,106 ,4 ,2 ,75 ,75 ,107 ,107 ,4 ,2 ,76 ,76 ,108 ,108 ,4 ,2 ,77 ,77 ,109 ,109 ,4 ,2 ,78 ,78 ,110 ,110 ,4 ,2 ,79 ,79 ,111 ,111 ,4 ,2 ,80 ,80 ,112 ,112 ,4 ,2 ,81 ,81 ,113 ,113 ,4 ,2 ,82 ,82 ,114 ,114 ,4 ,2 ,83 ,83 ,115 ,115 ,4 ,2 ,84 ,84 ,116 ,116 ,4 ,2 ,85 ,85 ,117 ,117 ,4 ,2 ,86 ,86 ,118 ,118 ,4 ,2 ,87 ,87 ,119 ,119 ,4 ,2 ,88 ,88 ,120 ,120 ,4 ,2 ,89 ,89 ,121 ,121 ,4 ,2 ,90 ,90 ,122 ,122 ,4 ,2 ,91 ,91 ,123 ,123 ,4 ,2 ,92 ,92 ,124 ,124 ,2 ,996 ,2 ,3 ,3 ,2 ,2 ,2 ,2 ,5 ,3 ,2 ,2 ,2 ,2 ,7 ,3 ,2 ,2 ,2 ,2 ,9 ,3 ,2 ,2 ,2 ,2 ,11 ,3 ,2 ,2 ,2 ,2 ,13 ,3 ,2 ,2 ,2 ,2 ,15 ,3 ,2 ,2 ,2 ,2 ,17 ,3 ,2 ,2 ,2 ,2 ,19 ,3 ,2 ,2 ,2 ,2 ,21 ,3 ,2 ,2 ,2 ,2 ,23 ,3 ,2 ,2 ,2 ,2 ,25 ,3 ,2 ,2 ,2 ,2 ,27 ,3 ,2 ,2 ,2 ,2 ,29 ,3 ,2 ,2 ,2 ,2 ,31 ,3 ,2 ,2 ,2 ,2 ,33 ,3 ,2 ,2 ,2 ,2 ,35 ,3 ,2 ,2 ,2 ,2 ,37 ,3 ,2 ,2 ,2 ,2 ,39 ,3 ,2 ,2 ,2 ,2 ,41 ,3 ,2 ,2 ,2 ,2 ,43 ,3 ,2 ,2 ,2 ,2 ,45 ,3 ,2 ,2 ,2 ,2 ,47 ,3 ,2 ,2 ,2 ,2 ,49 ,3 ,2 ,2 ,2 ,2 ,51 ,3 ,2 ,2 ,2 ,2 ,53 ,3 ,2 ,2 ,2 ,2 ,55 ,3 ,2 ,2 ,2 ,2 ,57 ,3 ,2 ,2 ,2 ,2 ,59 ,3 ,2 ,2 ,2 ,2 ,61 ,3 ,2 ,2 ,2 ,2 ,63 ,3 ,2 ,2 ,2 ,2 ,65 ,3 ,2 ,2 ,2 ,2 ,67 ,3 ,2 ,2 ,2 ,2 ,69 ,3 ,2 ,2 ,2 ,2 ,71 ,3 ,2 ,2 ,2 ,2 ,73 ,3 ,2 ,2 ,2 ,2 ,75 ,3 ,2 ,2 ,2 ,2 ,77 ,3 ,2 ,2 ,2 ,2 ,79 ,3 ,2 ,2 ,2 ,2 ,81 ,3 ,2 ,2 ,2 ,2 ,83 ,3 ,2 ,2 ,2 ,2 ,85 ,3 ,2 ,2 ,2 ,2 ,87 ,3 ,2 ,2 ,2 ,2 ,89 ,3 ,2 ,2 ,2 ,2 ,91 ,3 ,2 ,2 ,2 ,2 ,93 ,3 ,2 ,2 ,2 ,2 ,95 ,3 ,2 ,2 ,2 ,2 ,97 ,3 ,2 ,2 ,2 ,2 ,99 ,3 ,2 ,2 ,2 ,2 ,101 ,3 ,2 ,2 ,2 ,2 ,103 ,3 ,2 ,2 ,2 ,2 ,105 ,3 ,2 ,2 ,2 ,2 ,107 ,3 ,2 ,2 ,2 ,2 ,109 ,3 ,2 ,2 ,2 ,2 ,111 ,3 ,2 ,2 ,2 ,2 ,113 ,3 ,2 ,2 ,2 ,2 ,115 ,3 ,2 ,2 ,2 ,2 ,117 ,3 ,2 ,2 ,2 ,2 ,119 ,3 ,2 ,2 ,2 ,2 ,121 ,3 ,2 ,2 ,2 ,2 ,123 ,3 ,2 ,2 ,2 ,2 ,125 ,3 ,2 ,2 ,2 ,2 ,127 ,3 ,2 ,2 ,2 ,2 ,129 ,3 ,2 ,2 ,2 ,2 ,131 ,3 ,2 ,2 ,2 ,2 ,133 ,3 ,2 ,2 ,2 ,2 ,135 ,3 ,2 ,2 ,2 ,2 ,137 ,3 ,2 ,2 ,2 ,2 ,139 ,3 ,2 ,2 ,2 ,2 ,141 ,3 ,2 ,2 ,2 ,2 ,143 ,3 ,2 ,2 ,2 ,2 ,145 ,3 ,2 ,2 ,2 ,2 ,147 ,3 ,2 ,2 ,2 ,2 ,149 ,3 ,2 ,2 ,2 ,2 ,151 ,3 ,2 ,2 ,2 ,2 ,153 ,3 ,2 ,2 ,2 ,2 ,155 ,3 ,2 ,2 ,2 ,2 ,157 ,3 ,2 ,2 ,2 ,2 ,159 ,3 ,2 ,2 ,2 ,2 ,161 ,3 ,2 ,2 ,2 ,2 ,163 ,3 ,2 ,2 ,2 ,2 ,165 ,3 ,2 ,2 ,2 ,2 ,167 ,3 ,2 ,2 ,2 ,2 ,169 ,3 ,2 ,2 ,2 ,2 ,171 ,3 ,2 ,2 ,2 ,2 ,173 ,3 ,2 ,2 ,2 ,2 ,175 ,3 ,2 ,2 ,2 ,2 ,177 ,3 ,2 ,2 ,2 ,2 ,179 ,3 ,2 ,2 ,2 ,2 ,181 ,3 ,2 ,2 ,2 ,2 ,183 ,3 ,2 ,2 ,2 ,2 ,185 ,3 ,2 ,2 ,2 ,2 ,187 ,3 ,2 ,2 ,2 ,2 ,189 ,3 ,2 ,2 ,2 ,2 ,191 ,3 ,2 ,2 ,2 ,2 ,193 ,3 ,2 ,2 ,2 ,2 ,195 ,3 ,2 ,2 ,2 ,2 ,197 ,3 ,2 ,2 ,2 ,3 ,259 ,3 ,2 ,2 ,2 ,5 ,261 ,3 ,2 ,2 ,2 ,7 ,263 ,3 ,2 ,2 ,2 ,9 ,265 ,3 ,2 ,2 ,2 ,11 ,267 ,3 ,2 ,2 ,2 ,13 ,269 ,3 ,2 ,2 ,2 ,15 ,271 ,3 ,2 ,2 ,2 ,17 ,273 ,3 ,2 ,2 ,2 ,19 ,275 ,3 ,2 ,2 ,2 ,21 ,279 ,3 ,2 ,2 ,2 ,23 ,281 ,3 ,2 ,2 ,2 ,25 ,284 ,3 ,2 ,2 ,2 ,27 ,286 ,3 ,2 ,2 ,2 ,29 ,289 ,3 ,2 ,2 ,2 ,31 ,291 ,3 ,2 ,2 ,2 ,33 ,294 ,3 ,2 ,2 ,2 ,35 ,297 ,3 ,2 ,2 ,2 ,37 ,301 ,3 ,2 ,2 ,2 ,39 ,304 ,3 ,2 ,2 ,2 ,41 ,307 ,3 ,2 ,2 ,2 ,43 ,310 ,3 ,2 ,2 ,2 ,45 ,313 ,3 ,2 ,2 ,2 ,47 ,316 ,3 ,2 ,2 ,2 ,49 ,318 ,3 ,2 ,2 ,2 ,51 ,320 ,3 ,2 ,2 ,2 ,53 ,322 ,3 ,2 ,2 ,2 ,55 ,324 ,3 ,2 ,2 ,2 ,57 ,326 ,3 ,2 ,2 ,2 ,59 ,328 ,3 ,2 ,2 ,2 ,61 ,332 ,3 ,2 ,2 ,2 ,63 ,336 ,3 ,2 ,2 ,2 ,65 ,340 ,3 ,2 ,2 ,2 ,67 ,347 ,3 ,2 ,2 ,2 ,69 ,350 ,3 ,2 ,2 ,2 ,71 ,358 ,3 ,2 ,2 ,2 ,73 ,367 ,3 ,2 ,2 ,2 ,75 ,375 ,3 ,2 ,2 ,2 ,77 ,384 ,3 ,2 ,2 ,2 ,79 ,392 ,3 ,2 ,2 ,2 ,81 ,401 ,3 ,2 ,2 ,2 ,83 ,410 ,3 ,2 ,2 ,2 ,85 ,415 ,3 ,2 ,2 ,2 ,87 ,424 ,3 ,2 ,2 ,2 ,89 ,431 ,3 ,2 ,2 ,2 ,91 ,437 ,3 ,2 ,2 ,2 ,93 ,441 ,3 ,2 ,2 ,2 ,95 ,444 ,3 ,2 ,2 ,2 ,97 ,452 ,3 ,2 ,2 ,2 ,99 ,455 ,3 ,2 ,2 ,2 ,101 ,462 ,3 ,2 ,2 ,2 ,103 ,472 ,3 ,2 ,2 ,2 ,105 ,479 ,3 ,2 ,2 ,2 ,107 ,486 ,3 ,2 ,2 ,2 ,109 ,496 ,3 ,2 ,2 ,2 ,111 ,508 ,3 ,2 ,2 ,2 ,113 ,512 ,3 ,2 ,2 ,2 ,115 ,517 ,3 ,2 ,2 ,2 ,117 ,523 ,3 ,2 ,2 ,2 ,119 ,529 ,3 ,2 ,2 ,2 ,121 ,535 ,3 ,2 ,2 ,2 ,123 ,539 ,3 ,2 ,2 ,2 ,125 ,543 ,3 ,2 ,2 ,2 ,127 ,554 ,3 ,2 ,2 ,2 ,129 ,559 ,3 ,2 ,2 ,2 ,131 ,562 ,3 ,2 ,2 ,2 ,133 ,568 ,3 ,2 ,2 ,2 ,135 ,574 ,3 ,2 ,2 ,2 ,137 ,585 ,3 ,2 ,2 ,2 ,139 ,594 ,3 ,2 ,2 ,2 ,141 ,602 ,3 ,2 ,2 ,2 ,143 ,610 ,3 ,2 ,2 ,2 ,145 ,616 ,3 ,2 ,2 ,2 ,147 ,621 ,3 ,2 ,2 ,2 ,149 ,627 ,3 ,2 ,2 ,2 ,151 ,638 ,3 ,2 ,2 ,2 ,153 ,647 ,3 ,2 ,2 ,2 ,155 ,654 ,3 ,2 ,2 ,2 ,157 ,661 ,3 ,2 ,2 ,2 ,159 ,665 ,3 ,2 ,2 ,2 ,161 ,670 ,3 ,2 ,2 ,2 ,163 ,679 ,3 ,2 ,2 ,2 ,165 ,689 ,3 ,2 ,2 ,2 ,167 ,695 ,3 ,2 ,2 ,2 ,169 ,702 ,3 ,2 ,2 ,2 ,171 ,708 ,3 ,2 ,2 ,2 ,173 ,723 ,3 ,2 ,2 ,2 ,175 ,746 ,3 ,2 ,2 ,2 ,177 ,760 ,3 ,2 ,2 ,2 ,179 ,804 ,3 ,2 ,2 ,2 ,181 ,815 ,3 ,2 ,2 ,2 ,183 ,818 ,3 ,2 ,2 ,2 ,185 ,828 ,3 ,2 ,2 ,2 ,187 ,836 ,3 ,2 ,2 ,2 ,189 ,847 ,3 ,2 ,2 ,2 ,191 ,855 ,3 ,2 ,2 ,2 ,193 ,866 ,3 ,2 ,2 ,2 ,195 ,882 ,3 ,2 ,2 ,2 ,197 ,886 ,3 ,2 ,2 ,2 ,199 ,888 ,3 ,2 ,2 ,2 ,201 ,890 ,3 ,2 ,2 ,2 ,203 ,893 ,3 ,2 ,2 ,2 ,205 ,895 ,3 ,2 ,2 ,2 ,207 ,940 ,3 ,2 ,2 ,2 ,209 ,942 ,3 ,2 ,2 ,2 ,211 ,944 ,3 ,2 ,2 ,2 ,213 ,946 ,3 ,2 ,2 ,2 ,215 ,948 ,3 ,2 ,2 ,2 ,217 ,950 ,3 ,2 ,2 ,2 ,219 ,952 ,3 ,2 ,2 ,2 ,221 ,954 ,3 ,2 ,2 ,2 ,223 ,956 ,3 ,2 ,2 ,2 ,225 ,958 ,3 ,2 ,2 ,2 ,227 ,960 ,3 ,2 ,2 ,2 ,229 ,962 ,3 ,2 ,2 ,2 ,231 ,964 ,3 ,2 ,2 ,2 ,233 ,966 ,3 ,2 ,2 ,2 ,235 ,968 ,3 ,2 ,2 ,2 ,237 ,970 ,3 ,2 ,2 ,2 ,239 ,972 ,3 ,2 ,2 ,2 ,241 ,974 ,3 ,2 ,2 ,2 ,243 ,976 ,3 ,2 ,2 ,2 ,245 ,978 ,3 ,2 ,2 ,2 ,247 ,980 ,3 ,2 ,2 ,2 ,249 ,982 ,3 ,2 ,2 ,2 ,251 ,984 ,3 ,2 ,2 ,2 ,253 ,986 ,3 ,2 ,2 ,2 ,255 ,988 ,3 ,2 ,2 ,2 ,257 ,990 ,3 ,2 ,2 ,2 ,259 ,260 ,7 ,61 ,2 ,2 ,260 ,4 ,3 ,2 ,2 ,2 ,261 ,262 ,7 ,46 ,2 ,2 ,262 ,6 ,3 ,2 ,2 ,2 ,263 ,264 ,7 ,47 ,2 ,2 ,264 ,8 ,3 ,2 ,2 ,2 ,265 ,266 ,7 ,45 ,2 ,2 ,266 ,10 ,3 ,2 ,2 ,2 ,267 ,268 ,7 ,42 ,2 ,2 ,268 ,12 ,3 ,2 ,2 ,2 ,269 ,270 ,7 ,43 ,2 ,2 ,270 ,14 ,3 ,2 ,2 ,2 ,271 ,272 ,7 ,35 ,2 ,2 ,272 ,16 ,3 ,2 ,2 ,2 ,273 ,274 ,7 ,128 ,2 ,2 ,274 ,18 ,3 ,2 ,2 ,2 ,275 ,276 ,7 ,63 ,2 ,2 ,276 ,277 ,7 ,63 ,2 ,2 ,277 ,278 ,7 ,63 ,2 ,2 ,278 ,20 ,3 ,2 ,2 ,2 ,279 ,280 ,7 ,62 ,2 ,2 ,280 ,22 ,3 ,2 ,2 ,2 ,281 ,282 ,7 ,62 ,2 ,2 ,282 ,283 ,7 ,63 ,2 ,2 ,283 ,24 ,3 ,2 ,2 ,2 ,284 ,285 ,7 ,64 ,2 ,2 ,285 ,26 ,3 ,2 ,2 ,2 ,286 ,287 ,7 ,64 ,2 ,2 ,287 ,288 ,7 ,63 ,2 ,2 ,288 ,28 ,3 ,2 ,2 ,2 ,289 ,290 ,7 ,63 ,2 ,2 ,290 ,30 ,3 ,2 ,2 ,2 ,291 ,292 ,7 ,63 ,2 ,2 ,292 ,293 ,7 ,63 ,2 ,2 ,293 ,32 ,3 ,2 ,2 ,2 ,294 ,295 ,7 ,35 ,2 ,2 ,295 ,296 ,7 ,63 ,2 ,2 ,296 ,34 ,3 ,2 ,2 ,2 ,297 ,298 ,7 ,35 ,2 ,2 ,298 ,299 ,7 ,63 ,2 ,2 ,299 ,300 ,7 ,63 ,2 ,2 ,300 ,36 ,3 ,2 ,2 ,2 ,301 ,302 ,7 ,62 ,2 ,2 ,302 ,303 ,7 ,64 ,2 ,2 ,303 ,38 ,3 ,2 ,2 ,2 ,304 ,305 ,7 ,40 ,2 ,2 ,305 ,306 ,7 ,40 ,2 ,2 ,306 ,40 ,3 ,2 ,2 ,2 ,307 ,308 ,7 ,126 ,2 ,2 ,308 ,309 ,7 ,126 ,2 ,2 ,309 ,42 ,3 ,2 ,2 ,2 ,310 ,311 ,7 ,62 ,2 ,2 ,311 ,312 ,7 ,62 ,2 ,2 ,312 ,44 ,3 ,2 ,2 ,2 ,313 ,314 ,7 ,64 ,2 ,2 ,314 ,315 ,7 ,64 ,2 ,2 ,315 ,46 ,3 ,2 ,2 ,2 ,316 ,317 ,7 ,40 ,2 ,2 ,317 ,48 ,3 ,2 ,2 ,2 ,318 ,319 ,7 ,126 ,2 ,2 ,319 ,50 ,3 ,2 ,2 ,2 ,320 ,321 ,7 ,96 ,2 ,2 ,321 ,52 ,3 ,2 ,2 ,2 ,322 ,323 ,7 ,44 ,2 ,2 ,323 ,54 ,3 ,2 ,2 ,2 ,324 ,325 ,7 ,49 ,2 ,2 ,325 ,56 ,3 ,2 ,2 ,2 ,326 ,327 ,7 ,39 ,2 ,2 ,327 ,58 ,3 ,2 ,2 ,2 ,328 ,329 ,5 ,207 ,104 ,2 ,329 ,330 ,5 ,209 ,105 ,2 ,330 ,331 ,5 ,243 ,122 ,2 ,331 ,60 ,3 ,2 ,2 ,2 ,332 ,333 ,5 ,207 ,104 ,2 ,333 ,334 ,5 ,233 ,117 ,2 ,334 ,335 ,5 ,213 ,107 ,2 ,335 ,62 ,3 ,2 ,2 ,2 ,336 ,337 ,5 ,207 ,104 ,2 ,337 ,338 ,5 ,243 ,122 ,2 ,338 ,339 ,5 ,211 ,106 ,2 ,339 ,64 ,3 ,2 ,2 ,2 ,340 ,341 ,5 ,209 ,105 ,2 ,341 ,342 ,5 ,223 ,112 ,2 ,342 ,343 ,5 ,233 ,117 ,2 ,343 ,344 ,5 ,207 ,104 ,2 ,344 ,345 ,5 ,241 ,121 ,2 ,345 ,346 ,5 ,255 ,128 ,2 ,346 ,66 ,3 ,2 ,2 ,2 ,347 ,348 ,5 ,209 ,105 ,2 ,348 ,349 ,5 ,255 ,128 ,2 ,349 ,68 ,3 ,2 ,2 ,2 ,350 ,351 ,5 ,211 ,106 ,2 ,351 ,352 ,5 ,215 ,108 ,2 ,352 ,353 ,5 ,223 ,112 ,2 ,353 ,354 ,5 ,229 ,115 ,2 ,354 ,355 ,5 ,223 ,112 ,2 ,355 ,356 ,5 ,233 ,117 ,2 ,356 ,357 ,5 ,219 ,110 ,2 ,357 ,70 ,3 ,2 ,2 ,2 ,358 ,359 ,5 ,211 ,106 ,2 ,359 ,360 ,5 ,235 ,118 ,2 ,360 ,361 ,5 ,207 ,104 ,2 ,361 ,362 ,5 ,229 ,115 ,2 ,362 ,363 ,5 ,215 ,108 ,2 ,363 ,364 ,5 ,243 ,122 ,2 ,364 ,365 ,5 ,211 ,106 ,2 ,365 ,366 ,5 ,215 ,108 ,2 ,366 ,72 ,3 ,2 ,2 ,2 ,367 ,368 ,5 ,211 ,106 ,2 ,368 ,369 ,5 ,235 ,118 ,2 ,369 ,370 ,5 ,233 ,117 ,2 ,370 ,371 ,5 ,249 ,125 ,2 ,371 ,372 ,5 ,215 ,108 ,2 ,372 ,373 ,5 ,241 ,121 ,2 ,373 ,374 ,5 ,245 ,123 ,2 ,374 ,74 ,3 ,2 ,2 ,2 ,375 ,376 ,5 ,211 ,106 ,2 ,376 ,377 ,5 ,235 ,118 ,2 ,377 ,378 ,5 ,233 ,117 ,2 ,378 ,379 ,5 ,245 ,123 ,2 ,379 ,380 ,5 ,207 ,104 ,2 ,380 ,381 ,5 ,223 ,112 ,2 ,381 ,382 ,5 ,233 ,117 ,2 ,382 ,383 ,5 ,243 ,122 ,2 ,383 ,76 ,3 ,2 ,2 ,2 ,384 ,385 ,5 ,213 ,107 ,2 ,385 ,386 ,5 ,207 ,104 ,2 ,386 ,387 ,5 ,245 ,123 ,2 ,387 ,388 ,5 ,215 ,108 ,2 ,388 ,389 ,5 ,207 ,104 ,2 ,389 ,390 ,5 ,213 ,107 ,2 ,390 ,391 ,5 ,213 ,107 ,2 ,391 ,78 ,3 ,2 ,2 ,2 ,392 ,393 ,5 ,213 ,107 ,2 ,393 ,394 ,5 ,207 ,104 ,2 ,394 ,395 ,5 ,245 ,123 ,2 ,395 ,396 ,5 ,215 ,108 ,2 ,396 ,397 ,5 ,213 ,107 ,2 ,397 ,398 ,5 ,223 ,112 ,2 ,398 ,399 ,5 ,217 ,109 ,2 ,399 ,400 ,5 ,217 ,109 ,2 ,400 ,80 ,3 ,2 ,2 ,2 ,401 ,402 ,5 ,213 ,107 ,2 ,402 ,403 ,5 ,207 ,104 ,2 ,403 ,404 ,5 ,245 ,123 ,2 ,404 ,405 ,5 ,215 ,108 ,2 ,405 ,406 ,5 ,237 ,119 ,2 ,406 ,407 ,5 ,207 ,104 ,2 ,407 ,408 ,5 ,241 ,121 ,2 ,408 ,409 ,5 ,245 ,123 ,2 ,409 ,82 ,3 ,2 ,2 ,2 ,410 ,411 ,5 ,213 ,107 ,2 ,411 ,412 ,5 ,215 ,108 ,2 ,412 ,413 ,5 ,243 ,122 ,2 ,413 ,414 ,5 ,211 ,106 ,2 ,414 ,84 ,3 ,2 ,2 ,2 ,415 ,416 ,5 ,215 ,108 ,2 ,416 ,417 ,5 ,233 ,117 ,2 ,417 ,418 ,5 ,213 ,107 ,2 ,418 ,419 ,5 ,243 ,122 ,2 ,419 ,420 ,5 ,251 ,126 ,2 ,420 ,421 ,5 ,223 ,112 ,2 ,421 ,422 ,5 ,245 ,123 ,2 ,422 ,423 ,5 ,221 ,111 ,2 ,423 ,86 ,3 ,2 ,2 ,2 ,424 ,425 ,5 ,217 ,109 ,2 ,425 ,426 ,5 ,223 ,112 ,2 ,426 ,427 ,5 ,229 ,115 ,2 ,427 ,428 ,5 ,245 ,123 ,2 ,428 ,429 ,5 ,215 ,108 ,2 ,429 ,430 ,5 ,241 ,121 ,2 ,430 ,88 ,3 ,2 ,2 ,2 ,431 ,432 ,5 ,217 ,109 ,2 ,432 ,433 ,5 ,229 ,115 ,2 ,433 ,434 ,5 ,235 ,118 ,2 ,434 ,435 ,5 ,235 ,118 ,2 ,435 ,436 ,5 ,241 ,121 ,2 ,436 ,90 ,3 ,2 ,2 ,2 ,437 ,438 ,5 ,223 ,112 ,2 ,438 ,439 ,5 ,223 ,112 ,2 ,439 ,440 ,5 ,217 ,109 ,2 ,440 ,92 ,3 ,2 ,2 ,2 ,441 ,442 ,5 ,223 ,112 ,2 ,442 ,443 ,5 ,233 ,117 ,2 ,443 ,94 ,3 ,2 ,2 ,2 ,444 ,445 ,5 ,223 ,112 ,2 ,445 ,446 ,5 ,233 ,117 ,2 ,446 ,447 ,5 ,213 ,107 ,2 ,447 ,448 ,5 ,215 ,108 ,2 ,448 ,449 ,5 ,253 ,127 ,2 ,449 ,450 ,5 ,235 ,118 ,2 ,450 ,451 ,5 ,217 ,109 ,2 ,451 ,96 ,3 ,2 ,2 ,2 ,452 ,453 ,5 ,223 ,112 ,2 ,453 ,454 ,5 ,243 ,122 ,2 ,454 ,98 ,3 ,2 ,2 ,2 ,455 ,456 ,5 ,223 ,112 ,2 ,456 ,457 ,5 ,243 ,122 ,2 ,457 ,458 ,5 ,213 ,107 ,2 ,458 ,459 ,5 ,207 ,104 ,2 ,459 ,460 ,5 ,245 ,123 ,2 ,460 ,461 ,5 ,215 ,108 ,2 ,461 ,100 ,3 ,2 ,2 ,2 ,462 ,463 ,5 ,223 ,112 ,2 ,463 ,464 ,5 ,243 ,122 ,2 ,464 ,465 ,5 ,223 ,112 ,2 ,465 ,466 ,5 ,233 ,117 ,2 ,466 ,467 ,5 ,245 ,123 ,2 ,467 ,468 ,5 ,215 ,108 ,2 ,468 ,469 ,5 ,219 ,110 ,2 ,469 ,470 ,5 ,215 ,108 ,2 ,470 ,471 ,5 ,241 ,121 ,2 ,471 ,102 ,3 ,2 ,2 ,2 ,472 ,473 ,5 ,223 ,112 ,2 ,473 ,474 ,5 ,243 ,122 ,2 ,474 ,475 ,5 ,219 ,110 ,2 ,475 ,476 ,5 ,247 ,124 ,2 ,476 ,477 ,5 ,223 ,112 ,2 ,477 ,478 ,5 ,213 ,107 ,2 ,478 ,104 ,3 ,2 ,2 ,2 ,479 ,480 ,5 ,223 ,112 ,2 ,480 ,481 ,5 ,243 ,122 ,2 ,481 ,482 ,5 ,233 ,117 ,2 ,482 ,483 ,5 ,247 ,124 ,2 ,483 ,484 ,5 ,229 ,115 ,2 ,484 ,485 ,5 ,229 ,115 ,2 ,485 ,106 ,3 ,2 ,2 ,2 ,486 ,487 ,5 ,223 ,112 ,2 ,487 ,488 ,5 ,243 ,122 ,2 ,488 ,489 ,5 ,233 ,117 ,2 ,489 ,490 ,5 ,247 ,124 ,2 ,490 ,491 ,5 ,231 ,116 ,2 ,491 ,492 ,5 ,215 ,108 ,2 ,492 ,493 ,5 ,241 ,121 ,2 ,493 ,494 ,5 ,223 ,112 ,2 ,494 ,495 ,5 ,211 ,106 ,2 ,495 ,108 ,3 ,2 ,2 ,2 ,496 ,497 ,5 ,229 ,115 ,2 ,497 ,498 ,5 ,207 ,104 ,2 ,498 ,499 ,5 ,243 ,122 ,2 ,499 ,500 ,5 ,245 ,123 ,2 ,500 ,501 ,5 ,223 ,112 ,2 ,501 ,502 ,5 ,233 ,117 ,2 ,502 ,503 ,5 ,213 ,107 ,2 ,503 ,504 ,5 ,215 ,108 ,2 ,504 ,505 ,5 ,253 ,127 ,2 ,505 ,506 ,5 ,235 ,118 ,2 ,506 ,507 ,5 ,217 ,109 ,2 ,507 ,110 ,3 ,2 ,2 ,2 ,508 ,509 ,5 ,229 ,115 ,2 ,509 ,510 ,5 ,215 ,108 ,2 ,510 ,511 ,5 ,233 ,117 ,2 ,511 ,112 ,3 ,2 ,2 ,2 ,512 ,513 ,5 ,229 ,115 ,2 ,513 ,514 ,5 ,223 ,112 ,2 ,514 ,515 ,5 ,227 ,114 ,2 ,515 ,516 ,5 ,215 ,108 ,2 ,516 ,114 ,3 ,2 ,2 ,2 ,517 ,518 ,5 ,229 ,115 ,2 ,518 ,519 ,5 ,235 ,118 ,2 ,519 ,520 ,5 ,251 ,126 ,2 ,520 ,521 ,5 ,215 ,108 ,2 ,521 ,522 ,5 ,241 ,121 ,2 ,522 ,116 ,3 ,2 ,2 ,2 ,523 ,524 ,5 ,231 ,116 ,2 ,524 ,525 ,5 ,207 ,104 ,2 ,525 ,526 ,5 ,253 ,127 ,2 ,526 ,527 ,5 ,235 ,118 ,2 ,527 ,528 ,5 ,217 ,109 ,2 ,528 ,118 ,3 ,2 ,2 ,2 ,529 ,530 ,5 ,231 ,116 ,2 ,530 ,531 ,5 ,223 ,112 ,2 ,531 ,532 ,5 ,233 ,117 ,2 ,532 ,533 ,5 ,235 ,118 ,2 ,533 ,534 ,5 ,217 ,109 ,2 ,534 ,120 ,3 ,2 ,2 ,2 ,535 ,536 ,5 ,233 ,117 ,2 ,536 ,537 ,5 ,235 ,118 ,2 ,537 ,538 ,5 ,245 ,123 ,2 ,538 ,122 ,3 ,2 ,2 ,2 ,539 ,540 ,5 ,233 ,117 ,2 ,540 ,541 ,5 ,235 ,118 ,2 ,541 ,542 ,5 ,251 ,126 ,2 ,542 ,124 ,3 ,2 ,2 ,2 ,543 ,544 ,5 ,233 ,117 ,2 ,544 ,545 ,5 ,245 ,123 ,2 ,545 ,546 ,5 ,221 ,111 ,2 ,546 ,547 ,5 ,223 ,112 ,2 ,547 ,548 ,5 ,233 ,117 ,2 ,548 ,549 ,5 ,213 ,107 ,2 ,549 ,550 ,5 ,215 ,108 ,2 ,550 ,551 ,5 ,253 ,127 ,2 ,551 ,552 ,5 ,235 ,118 ,2 ,552 ,553 ,5 ,217 ,109 ,2 ,553 ,126 ,3 ,2 ,2 ,2 ,554 ,555 ,5 ,233 ,117 ,2 ,555 ,556 ,5 ,247 ,124 ,2 ,556 ,557 ,5 ,229 ,115 ,2 ,557 ,558 ,5 ,229 ,115 ,2 ,558 ,128 ,3 ,2 ,2 ,2 ,559 ,560 ,5 ,235 ,118 ,2 ,560 ,561 ,5 ,241 ,121 ,2 ,561 ,130 ,3 ,2 ,2 ,2 ,562 ,563 ,5 ,235 ,118 ,2 ,563 ,564 ,5 ,241 ,121 ,2 ,564 ,565 ,5 ,213 ,107 ,2 ,565 ,566 ,5 ,215 ,108 ,2 ,566 ,567 ,5 ,241 ,121 ,2 ,567 ,132 ,3 ,2 ,2 ,2 ,568 ,569 ,5 ,237 ,119 ,2 ,569 ,570 ,5 ,235 ,118 ,2 ,570 ,571 ,5 ,251 ,126 ,2 ,571 ,572 ,5 ,215 ,108 ,2 ,572 ,573 ,5 ,241 ,121 ,2 ,573 ,134 ,3 ,2 ,2 ,2 ,574 ,575 ,5 ,241 ,121 ,2 ,575 ,576 ,5 ,215 ,108 ,2 ,576 ,577 ,5 ,219 ,110 ,2 ,577 ,578 ,5 ,215 ,108 ,2 ,578 ,579 ,5 ,253 ,127 ,2 ,579 ,580 ,5 ,231 ,116 ,2 ,580 ,581 ,5 ,207 ,104 ,2 ,581 ,582 ,5 ,245 ,123 ,2 ,582 ,583 ,5 ,211 ,106 ,2 ,583 ,584 ,5 ,221 ,111 ,2 ,584 ,136 ,3 ,2 ,2 ,2 ,585 ,586 ,5 ,241 ,121 ,2 ,586 ,587 ,5 ,215 ,108 ,2 ,587 ,588 ,5 ,219 ,110 ,2 ,588 ,589 ,5 ,215 ,108 ,2 ,589 ,590 ,5 ,253 ,127 ,2 ,590 ,591 ,5 ,249 ,125 ,2 ,591 ,592 ,5 ,207 ,104 ,2 ,592 ,593 ,5 ,229 ,115 ,2 ,593 ,138 ,3 ,2 ,2 ,2 ,594 ,595 ,5 ,241 ,121 ,2 ,595 ,596 ,5 ,215 ,108 ,2 ,596 ,597 ,5 ,237 ,119 ,2 ,597 ,598 ,5 ,229 ,115 ,2 ,598 ,599 ,5 ,207 ,104 ,2 ,599 ,600 ,5 ,211 ,106 ,2 ,600 ,601 ,5 ,215 ,108 ,2 ,601 ,140 ,3 ,2 ,2 ,2 ,602 ,603 ,5 ,241 ,121 ,2 ,603 ,604 ,5 ,215 ,108 ,2 ,604 ,605 ,5 ,249 ,125 ,2 ,605 ,606 ,5 ,215 ,108 ,2 ,606 ,607 ,5 ,241 ,121 ,2 ,607 ,608 ,5 ,243 ,122 ,2 ,608 ,609 ,5 ,215 ,108 ,2 ,609 ,142 ,3 ,2 ,2 ,2 ,610 ,611 ,5 ,241 ,121 ,2 ,611 ,612 ,5 ,235 ,118 ,2 ,612 ,613 ,5 ,247 ,124 ,2 ,613 ,614 ,5 ,233 ,117 ,2 ,614 ,615 ,5 ,213 ,107 ,2 ,615 ,144 ,3 ,2 ,2 ,2 ,616 ,617 ,5 ,243 ,122 ,2 ,617 ,618 ,5 ,239 ,120 ,2 ,618 ,619 ,5 ,241 ,121 ,2 ,619 ,620 ,5 ,245 ,123 ,2 ,620 ,146 ,3 ,2 ,2 ,2 ,621 ,622 ,5 ,243 ,122 ,2 ,622 ,623 ,5 ,237 ,119 ,2 ,623 ,624 ,5 ,229 ,115 ,2 ,624 ,625 ,5 ,223 ,112 ,2 ,625 ,626 ,5 ,245 ,123 ,2 ,626 ,148 ,3 ,2 ,2 ,2 ,627 ,628 ,5 ,243 ,122 ,2 ,628 ,629 ,5 ,245 ,123 ,2 ,629 ,630 ,5 ,207 ,104 ,2 ,630 ,631 ,5 ,241 ,121 ,2 ,631 ,632 ,5 ,245 ,123 ,2 ,632 ,633 ,5 ,243 ,122 ,2 ,633 ,634 ,5 ,251 ,126 ,2 ,634 ,635 ,5 ,223 ,112 ,2 ,635 ,636 ,5 ,245 ,123 ,2 ,636 ,637 ,5 ,221 ,111 ,2 ,637 ,150 ,3 ,2 ,2 ,2 ,638 ,639 ,5 ,243 ,122 ,2 ,639 ,640 ,5 ,245 ,123 ,2 ,640 ,641 ,5 ,241 ,121 ,2 ,641 ,642 ,5 ,211 ,106 ,2 ,642 ,643 ,5 ,235 ,118 ,2 ,643 ,644 ,5 ,247 ,124 ,2 ,644 ,645 ,5 ,233 ,117 ,2 ,645 ,646 ,5 ,245 ,123 ,2 ,646 ,152 ,3 ,2 ,2 ,2 ,647 ,648 ,5 ,243 ,122 ,2 ,648 ,649 ,5 ,245 ,123 ,2 ,649 ,650 ,5 ,241 ,121 ,2 ,650 ,651 ,5 ,211 ,106 ,2 ,651 ,652 ,5 ,231 ,116 ,2 ,652 ,653 ,5 ,237 ,119 ,2 ,653 ,154 ,3 ,2 ,2 ,2 ,654 ,655 ,5 ,243 ,122 ,2 ,655 ,656 ,5 ,247 ,124 ,2 ,656 ,657 ,5 ,209 ,105 ,2 ,657 ,658 ,5 ,243 ,122 ,2 ,658 ,659 ,5 ,245 ,123 ,2 ,659 ,660 ,5 ,241 ,121 ,2 ,660 ,156 ,3 ,2 ,2 ,2 ,661 ,662 ,5 ,245 ,123 ,2 ,662 ,663 ,5 ,235 ,118 ,2 ,663 ,664 ,5 ,237 ,119 ,2 ,664 ,158 ,3 ,2 ,2 ,2 ,665 ,666 ,5 ,245 ,123 ,2 ,666 ,667 ,5 ,241 ,121 ,2 ,667 ,668 ,5 ,223 ,112 ,2 ,668 ,669 ,5 ,231 ,116 ,2 ,669 ,160 ,3 ,2 ,2 ,2 ,670 ,671 ,5 ,245 ,123 ,2 ,671 ,672 ,5 ,241 ,121 ,2 ,672 ,673 ,5 ,223 ,112 ,2 ,673 ,674 ,5 ,231 ,116 ,2 ,674 ,675 ,5 ,229 ,115 ,2 ,675 ,676 ,5 ,215 ,108 ,2 ,676 ,677 ,5 ,217 ,109 ,2 ,677 ,678 ,5 ,245 ,123 ,2 ,678 ,162 ,3 ,2 ,2 ,2 ,679 ,680 ,5 ,245 ,123 ,2 ,680 ,681 ,5 ,241 ,121 ,2 ,681 ,682 ,5 ,223 ,112 ,2 ,682 ,683 ,5 ,231 ,116 ,2 ,683 ,684 ,5 ,241 ,121 ,2 ,684 ,685 ,5 ,223 ,112 ,2 ,685 ,686 ,5 ,219 ,110 ,2 ,686 ,687 ,5 ,221 ,111 ,2 ,687 ,688 ,5 ,245 ,123 ,2 ,688 ,164 ,3 ,2 ,2 ,2 ,689 ,690 ,5 ,247 ,124 ,2 ,690 ,691 ,5 ,237 ,119 ,2 ,691 ,692 ,5 ,237 ,119 ,2 ,692 ,693 ,5 ,215 ,108 ,2 ,693 ,694 ,5 ,241 ,121 ,2 ,694 ,166 ,3 ,2 ,2 ,2 ,695 ,696 ,5 ,247 ,124 ,2 ,696 ,697 ,5 ,245 ,123 ,2 ,697 ,698 ,5 ,211 ,106 ,2 ,698 ,699 ,5 ,233 ,117 ,2 ,699 ,700 ,5 ,235 ,118 ,2 ,700 ,701 ,5 ,251 ,126 ,2 ,701 ,168 ,3 ,2 ,2 ,2 ,702 ,703 ,5 ,251 ,126 ,2 ,703 ,704 ,5 ,221 ,111 ,2 ,704 ,705 ,5 ,215 ,108 ,2 ,705 ,706 ,5 ,241 ,121 ,2 ,706 ,707 ,5 ,215 ,108 ,2 ,707 ,170 ,3 ,2 ,2 ,2 ,708 ,709 ,5 ,253 ,127 ,2 ,709 ,710 ,5 ,235 ,118 ,2 ,710 ,711 ,5 ,241 ,121 ,2 ,711 ,172 ,3 ,2 ,2 ,2 ,712 ,713 ,5 ,245 ,123 ,2 ,713 ,714 ,5 ,241 ,121 ,2 ,714 ,715 ,5 ,247 ,124 ,2 ,715 ,716 ,5 ,215 ,108 ,2 ,716 ,724 ,3 ,2 ,2 ,2 ,717 ,718 ,5 ,217 ,109 ,2 ,718 ,719 ,5 ,207 ,104 ,2 ,719 ,720 ,5 ,229 ,115 ,2 ,720 ,721 ,5 ,243 ,122 ,2 ,721 ,722 ,5 ,215 ,108 ,2 ,722 ,724 ,3 ,2 ,2 ,2 ,723 ,712 ,3 ,2 ,2 ,2 ,723 ,717 ,3 ,2 ,2 ,2 ,724 ,174 ,3 ,2 ,2 ,2 ,725 ,727 ,7 ,98 ,2 ,2 ,726 ,728 ,10 ,2 ,2 ,2 ,727 ,726 ,3 ,2 ,2 ,2 ,728 ,729 ,3 ,2 ,2 ,2 ,729 ,727 ,3 ,2 ,2 ,2 ,729 ,730 ,3 ,2 ,2 ,2 ,730 ,731 ,3 ,2 ,2 ,2 ,731 ,747 ,7 ,98 ,2 ,2 ,732 ,734 ,7 ,93 ,2 ,2 ,733 ,735 ,10 ,3 ,2 ,2 ,734 ,733 ,3 ,2 ,2 ,2 ,735 ,736 ,3 ,2 ,2 ,2 ,736 ,734 ,3 ,2 ,2 ,2 ,736 ,737 ,3 ,2 ,2 ,2 ,737 ,738 ,3 ,2 ,2 ,2 ,738 ,747 ,7 ,95 ,2 ,2 ,739 ,743 ,9 ,4 ,2 ,2 ,740 ,742 ,9 ,5 ,2 ,2 ,741 ,740 ,3 ,2 ,2 ,2 ,742 ,745 ,3 ,2 ,2 ,2 ,743 ,741 ,3 ,2 ,2 ,2 ,743 ,744 ,3 ,2 ,2 ,2 ,744 ,747 ,3 ,2 ,2 ,2 ,745 ,743 ,3 ,2 ,2 ,2 ,746 ,725 ,3 ,2 ,2 ,2 ,746 ,732 ,3 ,2 ,2 ,2 ,746 ,739 ,3 ,2 ,2 ,2 ,747 ,176 ,3 ,2 ,2 ,2 ,748 ,750 ,5 ,199 ,100 ,2 ,749 ,748 ,3 ,2 ,2 ,2 ,750 ,751 ,3 ,2 ,2 ,2 ,751 ,749 ,3 ,2 ,2 ,2 ,751 ,752 ,3 ,2 ,2 ,2 ,752 ,761 ,3 ,2 ,2 ,2 ,753 ,754 ,7 ,50 ,2 ,2 ,754 ,756 ,5 ,253 ,127 ,2 ,755 ,757 ,5 ,201 ,101 ,2 ,756 ,755 ,3 ,2 ,2 ,2 ,757 ,758 ,3 ,2 ,2 ,2 ,758 ,756 ,3 ,2 ,2 ,2 ,758 ,759 ,3 ,2 ,2 ,2 ,759 ,761 ,3 ,2 ,2 ,2 ,760 ,749 ,3 ,2 ,2 ,2 ,760 ,753 ,3 ,2 ,2 ,2 ,761 ,178 ,3 ,2 ,2 ,2 ,762 ,764 ,5 ,199 ,100 ,2 ,763 ,762 ,3 ,2 ,2 ,2 ,764 ,765 ,3 ,2 ,2 ,2 ,765 ,763 ,3 ,2 ,2 ,2 ,765 ,766 ,3 ,2 ,2 ,2 ,766 ,774 ,3 ,2 ,2 ,2 ,767 ,771 ,7 ,48 ,2 ,2 ,768 ,770 ,5 ,199 ,100 ,2 ,769 ,768 ,3 ,2 ,2 ,2 ,770 ,773 ,3 ,2 ,2 ,2 ,771 ,769 ,3 ,2 ,2 ,2 ,771 ,772 ,3 ,2 ,2 ,2 ,772 ,775 ,3 ,2 ,2 ,2 ,773 ,771 ,3 ,2 ,2 ,2 ,774 ,767 ,3 ,2 ,2 ,2 ,774 ,775 ,3 ,2 ,2 ,2 ,775 ,785 ,3 ,2 ,2 ,2 ,776 ,778 ,5 ,215 ,108 ,2 ,777 ,779 ,9 ,6 ,2 ,2 ,778 ,777 ,3 ,2 ,2 ,2 ,778 ,779 ,3 ,2 ,2 ,2 ,779 ,781 ,3 ,2 ,2 ,2 ,780 ,782 ,5 ,199 ,100 ,2 ,781 ,780 ,3 ,2 ,2 ,2 ,782 ,783 ,3 ,2 ,2 ,2 ,783 ,781 ,3 ,2 ,2 ,2 ,783 ,784 ,3 ,2 ,2 ,2 ,784 ,786 ,3 ,2 ,2 ,2 ,785 ,776 ,3 ,2 ,2 ,2 ,785 ,786 ,3 ,2 ,2 ,2 ,786 ,805 ,3 ,2 ,2 ,2 ,787 ,789 ,7 ,48 ,2 ,2 ,788 ,790 ,5 ,199 ,100 ,2 ,789 ,788 ,3 ,2 ,2 ,2 ,790 ,791 ,3 ,2 ,2 ,2 ,791 ,789 ,3 ,2 ,2 ,2 ,791 ,792 ,3 ,2 ,2 ,2 ,792 ,802 ,3 ,2 ,2 ,2 ,793 ,795 ,5 ,215 ,108 ,2 ,794 ,796 ,9 ,6 ,2 ,2 ,795 ,794 ,3 ,2 ,2 ,2 ,795 ,796 ,3 ,2 ,2 ,2 ,796 ,798 ,3 ,2 ,2 ,2 ,797 ,799 ,5 ,199 ,100 ,2 ,798 ,797 ,3 ,2 ,2 ,2 ,799 ,800 ,3 ,2 ,2 ,2 ,800 ,798 ,3 ,2 ,2 ,2 ,800 ,801 ,3 ,2 ,2 ,2 ,801 ,803 ,3 ,2 ,2 ,2 ,802 ,793 ,3 ,2 ,2 ,2 ,802 ,803 ,3 ,2 ,2 ,2 ,803 ,805 ,3 ,2 ,2 ,2 ,804 ,763 ,3 ,2 ,2 ,2 ,804 ,787 ,3 ,2 ,2 ,2 ,805 ,180 ,3 ,2 ,2 ,2 ,806 ,807 ,7 ,41 ,2 ,2 ,807 ,808 ,5 ,205 ,103 ,2 ,808 ,809 ,7 ,41 ,2 ,2 ,809 ,816 ,3 ,2 ,2 ,2 ,810 ,811 ,7 ,125 ,2 ,2 ,811 ,812 ,5 ,205 ,103 ,2 ,812 ,813 ,7 ,127 ,2 ,2 ,813 ,816 ,3 ,2 ,2 ,2 ,814 ,816 ,5 ,205 ,103 ,2 ,815 ,806 ,3 ,2 ,2 ,2 ,815 ,810 ,3 ,2 ,2 ,2 ,815 ,814 ,3 ,2 ,2 ,2 ,816 ,182 ,3 ,2 ,2 ,2 ,817 ,819 ,5 ,203 ,102 ,2 ,818 ,817 ,3 ,2 ,2 ,2 ,819 ,820 ,3 ,2 ,2 ,2 ,820 ,818 ,3 ,2 ,2 ,2 ,820 ,821 ,3 ,2 ,2 ,2 ,821 ,822 ,3 ,2 ,2 ,2 ,822 ,824 ,7 ,60 ,2 ,2 ,823 ,825 ,5 ,199 ,100 ,2 ,824 ,823 ,3 ,2 ,2 ,2 ,825 ,826 ,3 ,2 ,2 ,2 ,826 ,824 ,3 ,2 ,2 ,2 ,826 ,827 ,3 ,2 ,2 ,2 ,827 ,184 ,3 ,2 ,2 ,2 ,828 ,830 ,7 ,36 ,2 ,2 ,829 ,831 ,5 ,203 ,102 ,2 ,830 ,829 ,3 ,2 ,2 ,2 ,831 ,832 ,3 ,2 ,2 ,2 ,832 ,830 ,3 ,2 ,2 ,2 ,832 ,833 ,3 ,2 ,2 ,2 ,833 ,834 ,3 ,2 ,2 ,2 ,834 ,835 ,7 ,36 ,2 ,2 ,835 ,186 ,3 ,2 ,2 ,2 ,836 ,842 ,7 ,41 ,2 ,2 ,837 ,841 ,10 ,7 ,2 ,2 ,838 ,839 ,7 ,41 ,2 ,2 ,839 ,841 ,7 ,41 ,2 ,2 ,840 ,837 ,3 ,2 ,2 ,2 ,840 ,838 ,3 ,2 ,2 ,2 ,841 ,844 ,3 ,2 ,2 ,2 ,842 ,840 ,3 ,2 ,2 ,2 ,842 ,843 ,3 ,2 ,2 ,2 ,843 ,845 ,3 ,2 ,2 ,2 ,844 ,842 ,3 ,2 ,2 ,2 ,845 ,846 ,7 ,41 ,2 ,2 ,846 ,188 ,3 ,2 ,2 ,2 ,847 ,849 ,7 ,37 ,2 ,2 ,848 ,850 ,10 ,8 ,2 ,2 ,849 ,848 ,3 ,2 ,2 ,2 ,850 ,851 ,3 ,2 ,2 ,2 ,851 ,849 ,3 ,2 ,2 ,2 ,851 ,852 ,3 ,2 ,2 ,2 ,852 ,853 ,3 ,2 ,2 ,2 ,853 ,854 ,7 ,37 ,2 ,2 ,854 ,190 ,3 ,2 ,2 ,2 ,855 ,856 ,7 ,47 ,2 ,2 ,856 ,857 ,7 ,47 ,2 ,2 ,857 ,861 ,3 ,2 ,2 ,2 ,858 ,860 ,10 ,9 ,2 ,2 ,859 ,858 ,3 ,2 ,2 ,2 ,860 ,863 ,3 ,2 ,2 ,2 ,861 ,859 ,3 ,2 ,2 ,2 ,861 ,862 ,3 ,2 ,2 ,2 ,862 ,864 ,3 ,2 ,2 ,2 ,863 ,861 ,3 ,2 ,2 ,2 ,864 ,865 ,8 ,96 ,2 ,2 ,865 ,192 ,3 ,2 ,2 ,2 ,866 ,867 ,7 ,49 ,2 ,2 ,867 ,868 ,7 ,44 ,2 ,2 ,868 ,872 ,3 ,2 ,2 ,2 ,869 ,871 ,11 ,2 ,2 ,2 ,870 ,869 ,3 ,2 ,2 ,2 ,871 ,874 ,3 ,2 ,2 ,2 ,872 ,873 ,3 ,2 ,2 ,2 ,872 ,870 ,3 ,2 ,2 ,2 ,873 ,878 ,3 ,2 ,2 ,2 ,874 ,872 ,3 ,2 ,2 ,2 ,875 ,876 ,7 ,44 ,2 ,2 ,876 ,879 ,7 ,49 ,2 ,2 ,877 ,879 ,7 ,2 ,2 ,3 ,878 ,875 ,3 ,2 ,2 ,2 ,878 ,877 ,3 ,2 ,2 ,2 ,879 ,880 ,3 ,2 ,2 ,2 ,880 ,881 ,8 ,97 ,2 ,2 ,881 ,194 ,3 ,2 ,2 ,2 ,882 ,883 ,9 ,10 ,2 ,2 ,883 ,884 ,3 ,2 ,2 ,2 ,884 ,885 ,8 ,98 ,2 ,2 ,885 ,196 ,3 ,2 ,2 ,2 ,886 ,887 ,11 ,2 ,2 ,2 ,887 ,198 ,3 ,2 ,2 ,2 ,888 ,889 ,9 ,11 ,2 ,2 ,889 ,200 ,3 ,2 ,2 ,2 ,890 ,891 ,9 ,12 ,2 ,2 ,891 ,202 ,3 ,2 ,2 ,2 ,892 ,894 ,9 ,13 ,2 ,2 ,893 ,892 ,3 ,2 ,2 ,2 ,894 ,204 ,3 ,2 ,2 ,2 ,895 ,896 ,5 ,201 ,101 ,2 ,896 ,897 ,5 ,201 ,101 ,2 ,897 ,898 ,5 ,201 ,101 ,2 ,898 ,899 ,5 ,201 ,101 ,2 ,899 ,900 ,5 ,201 ,101 ,2 ,900 ,901 ,5 ,201 ,101 ,2 ,901 ,902 ,5 ,201 ,101 ,2 ,902 ,904 ,5 ,201 ,101 ,2 ,903 ,905 ,7 ,47 ,2 ,2 ,904 ,903 ,3 ,2 ,2 ,2 ,904 ,905 ,3 ,2 ,2 ,2 ,905 ,906 ,3 ,2 ,2 ,2 ,906 ,907 ,5 ,201 ,101 ,2 ,907 ,908 ,5 ,201 ,101 ,2 ,908 ,909 ,5 ,201 ,101 ,2 ,909 ,911 ,5 ,201 ,101 ,2 ,910 ,912 ,7 ,47 ,2 ,2 ,911 ,910 ,3 ,2 ,2 ,2 ,911 ,912 ,3 ,2 ,2 ,2 ,912 ,913 ,3 ,2 ,2 ,2 ,913 ,914 ,5 ,201 ,101 ,2 ,914 ,915 ,5 ,201 ,101 ,2 ,915 ,916 ,5 ,201 ,101 ,2 ,916 ,918 ,5 ,201 ,101 ,2 ,917 ,919 ,7 ,47 ,2 ,2 ,918 ,917 ,3 ,2 ,2 ,2 ,918 ,919 ,3 ,2 ,2 ,2 ,919 ,920 ,3 ,2 ,2 ,2 ,920 ,921 ,5 ,201 ,101 ,2 ,921 ,922 ,5 ,201 ,101 ,2 ,922 ,923 ,5 ,201 ,101 ,2 ,923 ,925 ,5 ,201 ,101 ,2 ,924 ,926 ,7 ,47 ,2 ,2 ,925 ,924 ,3 ,2 ,2 ,2 ,925 ,926 ,3 ,2 ,2 ,2 ,926 ,927 ,3 ,2 ,2 ,2 ,927 ,928 ,5 ,201 ,101 ,2 ,928 ,929 ,5 ,201 ,101 ,2 ,929 ,930 ,5 ,201 ,101 ,2 ,930 ,931 ,5 ,201 ,101 ,2 ,931 ,932 ,5 ,201 ,101 ,2 ,932 ,933 ,5 ,201 ,101 ,2 ,933 ,934 ,5 ,201 ,101 ,2 ,934 ,935 ,5 ,201 ,101 ,2 ,935 ,936 ,5 ,201 ,101 ,2 ,936 ,937 ,5 ,201 ,101 ,2 ,937 ,938 ,5 ,201 ,101 ,2 ,938 ,939 ,5 ,201 ,101 ,2 ,939 ,206 ,3 ,2 ,2 ,2 ,940 ,941 ,9 ,14 ,2 ,2 ,941 ,208 ,3 ,2 ,2 ,2 ,942 ,943 ,9 ,15 ,2 ,2 ,943 ,210 ,3 ,2 ,2 ,2 ,944 ,945 ,9 ,16 ,2 ,2 ,945 ,212 ,3 ,2 ,2 ,2 ,946 ,947 ,9 ,17 ,2 ,2 ,947 ,214 ,3 ,2 ,2 ,2 ,948 ,949 ,9 ,18 ,2 ,2 ,949 ,216 ,3 ,2 ,2 ,2 ,950 ,951 ,9 ,19 ,2 ,2 ,951 ,218 ,3 ,2 ,2 ,2 ,952 ,953 ,9 ,20 ,2 ,2 ,953 ,220 ,3 ,2 ,2 ,2 ,954 ,955 ,9 ,21 ,2 ,2 ,955 ,222 ,3 ,2 ,2 ,2 ,956 ,957 ,9 ,22 ,2 ,2 ,957 ,224 ,3 ,2 ,2 ,2 ,958 ,959 ,9 ,23 ,2 ,2 ,959 ,226 ,3 ,2 ,2 ,2 ,960 ,961 ,9 ,24 ,2 ,2 ,961 ,228 ,3 ,2 ,2 ,2 ,962 ,963 ,9 ,25 ,2 ,2 ,963 ,230 ,3 ,2 ,2 ,2 ,964 ,965 ,9 ,26 ,2 ,2 ,965 ,232 ,3 ,2 ,2 ,2 ,966 ,967 ,9 ,27 ,2 ,2 ,967 ,234 ,3 ,2 ,2 ,2 ,968 ,969 ,9 ,28 ,2 ,2 ,969 ,236 ,3 ,2 ,2 ,2 ,970 ,971 ,9 ,29 ,2 ,2 ,971 ,238 ,3 ,2 ,2 ,2 ,972 ,973 ,9 ,30 ,2 ,2 ,973 ,240 ,3 ,2 ,2 ,2 ,974 ,975 ,9 ,31 ,2 ,2 ,975 ,242 ,3 ,2 ,2 ,2 ,976 ,977 ,9 ,32 ,2 ,2 ,977 ,244 ,3 ,2 ,2 ,2 ,978 ,979 ,9 ,33 ,2 ,2 ,979 ,246 ,3 ,2 ,2 ,2 ,980 ,981 ,9 ,34 ,2 ,2 ,981 ,248 ,3 ,2 ,2 ,2 ,982 ,983 ,9 ,35 ,2 ,2 ,983 ,250 ,3 ,2 ,2 ,2 ,984 ,985 ,9 ,36 ,2 ,2 ,985 ,252 ,3 ,2 ,2 ,2 ,986 ,987 ,9 ,37 ,2 ,2 ,987 ,254 ,3 ,2 ,2 ,2 ,988 ,989 ,9 ,38 ,2 ,2 ,989 ,256 ,3 ,2 ,2 ,2 ,990 ,991 ,9 ,39 ,2 ,2 ,991 ,258 ,3 ,2 ,2 ,2 ,37 ,2 ,723 ,729 ,736 ,743 ,746 ,751 ,758 ,760 ,765 ,771 ,774 ,778 ,783 ,785 ,791 ,795 ,800 ,802 ,804 ,815 ,820 ,826 ,832 ,840 ,842 ,851 ,861 ,872 ,878 ,893 ,904 ,911 ,918 ,925 ,3 ,2 ,3 ,2 ] 
lexer_channel_names=["DEFAULT_TOKEN_CHANNEL" ,"HIDDEN" ] 
lexer_mode_names=["DEFAULT_MODE" ] 
lexer_literal_names=["" ,"';'" ,"','" ,"'-'" ,"'+'" ,"'('" ,"')'" ,"'!'" ,"'~'" ,"'==='" ,"'<'" ,"'<='" ,"'>'" ,"'>='" ,"'='" ,"'=='" ,"'!='" ,"'!=='" ,"'<>'" ,"'&&'" ,"'||'" ,"'<<'" ,"'>>'" ,"'&'" ,"'|'" ,"'^'" ,"'*'" ,"'/'" ,"'%'" ] 
lexer_symbolic_names=["" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"" ,"K_ABS" ,"K_AND" ,"K_ASC" ,"K_BINARY" ,"K_BY" ,"K_CEILING" ,"K_COALESCE" ,"K_CONVERT" ,"K_CONTAINS" ,"K_DATEADD" ,"K_DATEDIFF" ,"K_DATEPART" ,"K_DESC" ,"K_ENDSWITH" ,"K_FILTER" ,"K_FLOOR" ,"K_IIF" ,"K_IN" ,"K_INDEXOF" ,"K_IS" ,"K_ISDATE" ,"K_ISINTEGER" ,"K_ISGUID" ,"K_ISNULL" ,"K_ISNUMERIC" ,"K_LASTINDEXOF" ,"K_LEN" ,"K_LIKE" ,"K_LOWER" ,"K_MAXOF" ,"K_MINOF" ,"K_NOT" ,"K_NOW" ,"K_NTHINDEXOF" ,"K_NULL" ,"K_OR" ,"K_ORDER" ,"K_POWER" ,"K_REGEXMATCH" ,"K_REGEXVAL" ,"K_REPLACE" ,"K_REVERSE" ,"K_ROUND" ,"K_SQRT" ,"K_SPLIT" ,"K_STARTSWITH" ,"K_STRCOUNT" ,"K_STRCMP" ,"K_SUBSTR" ,"K_TOP" ,"K_TRIM" ,"K_TRIMLEFT" ,"K_TRIMRIGHT" ,"K_UPPER" ,"K_UTCNOW" ,"K_WHERE" ,"K_XOR" ,"BOOLEAN_LITERAL" ,"IDENTIFIER" ,"INTEGER_LITERAL" ,"NUMERIC_LITERAL" ,"GUID_LITERAL" ,"MEASUREMENT_KEY_LITERAL" ,"POINT_TAG_LITERAL" ,"STRING_LITERAL" ,"DATETIME_LITERAL" ,"SINGLE_LINE_COMMENT" ,"MULTILINE_COMMENT" ,"SPACES" ,"UNEXPECTED_CHAR" ] 
lexer_rule_names=["T__0" ,"T__1" ,"T__2" ,"T__3" ,"T__4" ,"T__5" ,"T__6" ,"T__7" ,"T__8" ,"T__9" ,"T__10" ,"T__11" ,"T__12" ,"T__13" ,"T__14" ,"T__15" ,"T__16" ,"T__17" ,"T__18" ,"T__19" ,"T__20" ,"T__21" ,"T__22" ,"T__23" ,"T__24" ,"T__25" ,"T__26" ,"T__27" ,"K_ABS" ,"K_AND" ,"K_ASC" ,"K_BINARY" ,"K_BY" ,"K_CEILING" ,"K_COALESCE" ,"K_CONVERT" ,"K_CONTAINS" ,"K_DATEADD" ,"K_DATEDIFF" ,"K_DATEPART" ,"K_DESC" ,"K_ENDSWITH" ,"K_FILTER" ,"K_FLOOR" ,"K_IIF" ,"K_IN" ,"K_INDEXOF" ,"K_IS" ,"K_ISDATE" ,"K_ISINTEGER" ,"K_ISGUID" ,"K_ISNULL" ,"K_ISNUMERIC" ,"K_LASTINDEXOF" ,"K_LEN" ,"K_LIKE" ,"K_LOWER" ,"K_MAXOF" ,"K_MINOF" ,"K_NOT" ,"K_NOW" ,"K_NTHINDEXOF" ,"K_NULL" ,"K_OR" ,"K_ORDER" ,"K_POWER" ,"K_REGEXMATCH" ,"K_REGEXVAL" ,"K_REPLACE" ,"K_REVERSE" ,"K_ROUND" ,"K_SQRT" ,"K_SPLIT" ,"K_STARTSWITH" ,"K_STRCOUNT" ,"K_STRCMP" ,"K_SUBSTR" ,"K_TOP" ,"K_TRIM" ,"K_TRIMLEFT" ,"K_TRIMRIGHT" ,"K_UPPER" ,"K_UTCNOW" ,"K_WHERE" ,"K_XOR" ,"BOOLEAN_LITERAL" ,"IDENTIFIER" ,"INTEGER_LITERAL" ,"NUMERIC_LITERAL" ,"GUID_LITERAL" ,"MEASUREMENT_KEY_LITERAL" ,"POINT_TAG_LITERAL" ,"STRING_LITERAL" ,"DATETIME_LITERAL" ,"SINGLE_LINE_COMMENT" ,"MULTILINE_COMMENT" ,"SPACES" ,"UNEXPECTED_CHAR" ,"DIGIT" ,"HEX_DIGIT" ,"ACRONYM_DIGIT" ,"GUID_VALUE" ,"A" ,"B" ,"C" ,"D" ,"E" ,"F" ,"G" ,"H" ,"I" ,"J" ,"K" ,"L" ,"M" ,"N" ,"O" ,"P" ,"Q" ,"R" ,"S" ,"T" ,"U" ,"V" ,"W" ,"X" ,"Y" ,"Z" ] 
filter_expression_syntax_lexer_t_0=1 
filter_expression_syntax_lexer_t_1=2 
filter_expression_syntax_lexer_t_2=3 
filter_expression_syntax_lexer_t_3=4 
filter_expression_syntax_lexer_t_4=5 
filter_expression_syntax_lexer_t_5=6 
filter_expression_syntax_lexer_t_6=7 
filter_expression_syntax_lexer_t_7=8 
filter_expression_syntax_lexer_t_8=9 
filter_expression_syntax_lexer_t_9=10 
filter_expression_syntax_lexer_t_10=11 
filter_expression_syntax_lexer_t_11=12 
filter_expression_syntax_lexer_t_12=13 
filter_expression_syntax_lexer_t_13=14 
filter_expression_syntax_lexer_t_14=15 
filter_expression_syntax_lexer_t_15=16 
filter_expression_syntax_lexer_t_16=17 
filter_expression_syntax_lexer_t_17=18 
filter_expression_syntax_lexer_t_18=19 
filter_expression_syntax_lexer_t_19=20 
filter_expression_syntax_lexer_t_20=21 
filter_expression_syntax_lexer_t_21=22 
filter_expression_syntax_lexer_t_22=23 
filter_expression_syntax_lexer_t_23=24 
filter_expression_syntax_lexer_t_24=25 
filter_expression_syntax_lexer_t_25=26 
filter_expression_syntax_lexer_t_26=27 
filter_expression_syntax_lexer_t_27=28 
filter_expression_syntax_lexer_k_abs=29 
filter_expression_syntax_lexer_k_and=30 
filter_expression_syntax_lexer_k_asc=31 
filter_expression_syntax_lexer_k_binary=32 
filter_expression_syntax_lexer_k_by=33 
filter_expression_syntax_lexer_k_ceiling=34 
filter_expression_syntax_lexer_k_coalesce=35 
filter_expression_syntax_lexer_k_convert=36 
filter_expression_syntax_lexer_k_contains=37 
filter_expression_syntax_lexer_k_dateadd=38 
filter_expression_syntax_lexer_k_datediff=39 
filter_expression_syntax_lexer_k_datepart=40 
filter_expression_syntax_lexer_k_desc=41 
filter_expression_syntax_lexer_k_endswith=42 
filter_expression_syntax_lexer_k_filter=43 
filter_expression_syntax_lexer_k_floor=44 
filter_expression_syntax_lexer_k_iif=45 
filter_expression_syntax_lexer_k_in=46 
filter_expression_syntax_lexer_k_indexof=47 
filter_expression_syntax_lexer_k_is=48 
filter_expression_syntax_lexer_k_isdate=49 
filter_expression_syntax_lexer_k_isinteger=50 
filter_expression_syntax_lexer_k_isguid=51 
filter_expression_syntax_lexer_k_isnull=52 
filter_expression_syntax_lexer_k_isnumeric=53 
filter_expression_syntax_lexer_k_lastindexof=54 
filter_expression_syntax_lexer_k_len=55 
filter_expression_syntax_lexer_k_like=56 
filter_expression_syntax_lexer_k_lower=57 
filter_expression_syntax_lexer_k_maxof=58 
filter_expression_syntax_lexer_k_minof=59 
filter_expression_syntax_lexer_k_not=60 
filter_expression_syntax_lexer_k_now=61 
filter_expression_syntax_lexer_k_nthindexof=62 
filter_expression_syntax_lexer_k_null=63 
filter_expression_syntax_lexer_k_or=64 
filter_expression_syntax_lexer_k_order=65 
filter_expression_syntax_lexer_k_power=66 
filter_expression_syntax_lexer_k_regexmatch=67 
filter_expression_syntax_lexer_k_regexval=68 
filter_expression_syntax_lexer_k_replace=69 
filter_expression_syntax_lexer_k_reverse=70 
filter_expression_syntax_lexer_k_round=71 
filter_expression_syntax_lexer_k_sqrt=72 
filter_expression_syntax_lexer_k_split=73 
filter_expression_syntax_lexer_k_startswith=74 
filter_expression_syntax_lexer_k_strcount=75 
filter_expression_syntax_lexer_k_strcmp=76 
filter_expression_syntax_lexer_k_substr=77 
filter_expression_syntax_lexer_k_top=78 
filter_expression_syntax_lexer_k_trim=79 
filter_expression_syntax_lexer_k_trimleft=80 
filter_expression_syntax_lexer_k_trimright=81 
filter_expression_syntax_lexer_k_upper=82 
filter_expression_syntax_lexer_k_utcnow=83 
filter_expression_syntax_lexer_k_where=84 
filter_expression_syntax_lexer_k_xor=85 
filter_expression_syntax_lexer_boolean_literal=86 
filter_expression_syntax_lexer_identifier=87 
filter_expression_syntax_lexer_integer_literal=88 
filter_expression_syntax_lexer_numeric_literal=89 
filter_expression_syntax_lexer_guid_literal=90 
filter_expression_syntax_lexer_measurement_key_literal=91 
filter_expression_syntax_lexer_point_tag_literal=92 
filter_expression_syntax_lexer_string_literal=93 
filter_expression_syntax_lexer_datetime_literal=94 
filter_expression_syntax_lexer_single_line_comment=95 
filter_expression_syntax_lexer_multiline_comment=96 
filter_expression_syntax_lexer_spaces=97 
filter_expression_syntax_lexer_unexpected_char=98 
)
struct FilterExpressionSyntaxLexer {&antlr.BaseLexer

mut:
channel_names []string 
mode_names []string 
}
// NewFilterExpressionSyntaxLexer produces a new lexer instance for the optional input antlr.CharStr
pub fn new_filter_expression_syntax_lexer(input antlr.CharStream) (&FilterExpressionSyntaxLexer, ) {mut l:=new(FilterExpressionSyntaxLexer ,)  
mut lexer_deserializer:=antlr.new_atndeserializer(unsafe { nil } ,)  
mut lexer_atn:=lexer_deserializer.deserialize_from_uint16(serialized_lexer_atn ,)  
mut lexer_decision_to_dfa:=[]*antlr.DFA{len: lexer_atn.decision_to_state .len }  
for index, ds in  lexer_atn.decision_to_state  {
lexer_decision_to_dfa[index ]=antlr.new_dfa(ds ,index ,)  
}
l.base_lexer=antlr.new_base_lexer(input ,)  
l.interpreter=antlr.new_lexer_atnsimulator(l ,lexer_atn ,lexer_decision_to_dfa ,antlr.new_prediction_context_cache() ,)  
l.channel_names=lexer_channel_names  
l.mode_names=lexer_mode_names  
l.rule_names=lexer_rule_names  
l.literal_names=lexer_literal_names  
l.symbolic_names=lexer_symbolic_names  
l.grammar_file_name="FilterExpressionSyntax.g4"  
return l 
}
