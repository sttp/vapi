module parser

import github.com.antlr.antlr4.runtime.Go.antlr
